-- Data Sampler (dataSampler.vhd)
-- Asynchronous reset, active high
------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.ALL;

ENTITY dataSampler IS
  PORT (
    clk: in STD_ULOGIC;
    reset: in STD_ULOGIC;
    outValid: out STD_ULOGIC;
    A_in: in STD_ULOGIC_VECTOR(7 DOWNTO 0);
    B_in: in STD_ULOGIC_VECTOR(7 DOWNTO 0);
    C_in: in STD_ULOGIC_VECTOR(7 DOWNTO 0);
    D_in: in STD_ULOGIC_VECTOR(7 DOWNTO 0);
    E_in: in STD_ULOGIC_VECTOR(7 DOWNTO 0);
    F_out: out STD_ULOGIC_VECTOR(15 DOWNTO 0);
    G_out: out STD_ULOGIC_VECTOR(15 DOWNTO 0)
  );
END;

ARCHITECTURE oneAdd_oneMult OF dataSampler IS
  TYPE MUXSEL is (LEFT, RIGHT);
  TYPE STATE_TYPE is (STAGE0, STAGE1, STAGE2, STAGE3, STAGE4);
  SIGNAL curState, nextState : STATE_TYPE;      
  -- control signals
  SIGNAL M1_sel, M2_sel, M3_sel : MUXSEL;
  SIGNAL R1_en, R2_en, R3_en, R4_en, R5_en, R6_en : BOOLEAN;
  -- data signals
  SIGNAL reg1_in, reg2_in, reg3_in: SIGNED(7 DOWNTO 0);
  SIGNAL reg1, reg2, reg3, reg4, addOut: SIGNED(7 DOWNTO 0);
  SIGNAL reg5, reg6, multOut : SIGNED(15 DOWNTO 0);
BEGIN
  
  M1: PROCESS(M1_sel,A_in,C_in)
  BEGIN
    IF M1_sel = LEFT THEN
      reg1_in <= signed(A_in);
    ELSE -- RIGHT
      reg1_in <= signed(C_in);
    END IF;
  END PROCESS;
  
  M2: PROCESS(M2_sel,B_in,D_in)
  BEGIN
    IF M2_sel = LEFT THEN
      reg2_in <= signed(B_in);
    ELSE -- RIGHT
      reg2_in <= signed(D_in);
    END IF;
  END PROCESS;
  
  M3: PROCESS(M3_sel,E_in,addOut)
  BEGIN
    IF M3_sel = LEFT THEN
      reg3_in <= signed(E_in);
    ELSE -- RIGHT
      reg3_in <= signed(addOut);
    END IF;
  END PROCESS;  
  
  R1: PROCESS(reset,clk)
  BEGIN
    IF reset = '1' THEN
      reg1 <= TO_SIGNED(0,8);
    ELSIF clk'event AND clk='1' THEN
      IF R1_en = true THEN
        reg1 <= reg1_in;
      END IF;
    END IF;
  END PROCESS;      
        
  R2: PROCESS(reset,clk)
  BEGIN
    IF reset = '1' THEN
      reg2 <= TO_SIGNED(0,8);
    ELSIF clk'event AND clk='1' THEN
      IF R2_en = true THEN
        reg2 <= reg2_in;
      END IF;
    END IF;
  END PROCESS;      
  
  R3: PROCESS(reset,clk)
  BEGIN
    IF reset = '1' THEN
      reg3 <= TO_SIGNED(0,8);
    ELSIF clk'event AND clk='1' THEN
      IF R3_en = true THEN --
        reg3 <= reg3_in;
      END IF;
    END IF;
  END PROCESS;      
        
  R4: PROCESS(reset,clk)
  BEGIN
    IF reset = '1' THEN
      reg4 <= TO_SIGNED(0,8);
    ELSIF clk'event AND clk='1' THEN
      IF R4_en = true THEN
        reg4 <= addOut;
      END IF;
    END IF;
  END PROCESS;

  add: PROCESS(reg1, reg2)
  BEGIN
    addOut <= reg1 + reg2;
  END PROCESS;        

  mult: PROCESS(reg3, reg4)
  BEGIN
    multOut <= reg3 * reg4;
  END PROCESS;        
  
  R5: PROCESS(reset,clk)
  BEGIN
    IF reset = '1' THEN
      reg5 <= TO_SIGNED(0,16);
    ELSIF clk'event and clk='1' THEN
      IF R5_en = true THEN
        reg5 <= multOut;
      END IF;
    END IF;
  END PROCESS;
  
  R6: PROCESS(reset,clk)
  BEGIN
    IF reset = '1' THEN
      reg6 <= TO_SIGNED(0,16);
    ELSIF clk'event AND clk='1' THEN
      IF R6_en = true THEN
        reg6 <= multOut;
      END IF;
    END IF;
  END PROCESS;

  F_out <= STD_ULOGIC_VECTOR(reg5); -- type casting
  G_out <= STD_ULOGIC_VECTOR(reg6);  
  
  stateReg: PROCESS(reset,clk)
  BEGIN
    IF reset = '1'  THEN
      curState <= STAGE0;
    ELSIF clk'event AND clk = '1' THEN
      curState <= nextState;
    END IF;
  END PROCESS;
  
  nextStateLogic: PROCESS(curState)
  BEGIN
    
    CASE curState IS
      WHEN STAGE0 =>
        if reg1 = reg1_in and reg2 = reg1_in then 
          nextState => STAGE1;
        else
          nextState => STAGE0;  
      end if; 
      WHEN STAGE1 =>
         if addOut = reg1 + reg2 then 
            nexState => STAGE2;
        else 
            reset = '1';
            nextState => STAGE0; 
     WHEN STAGE3 =>
       if reg3 = reg3_in and reg4 = addOut then 
          nextState => STAGE1;
     else
          nextState
    WHEN OTHERS => 
      nextState <= STAGE0;
    END CASE;
  END PROCESS;-- nextStateLogic
  
  ctrlOut: PROCESS(curState)
  BEGIN
    -- assign default values
    M1_sel <= ;
    M2_sel <= ;
    M3_sel <= ;
    
    R1_en, R2_en, R3_en, R4_en, R5_en, R6_en := FALSE ;

    outValid <= '0';
    CASE curState IS
      
      WHEN STAGE0 =>
        M1_sel = LEFT;
        M2_sel = LEFT;
      WHEN STAGE1 =>  
        M1_sel = RIGHT;
        M2_sel = RIGHT;
        M3_sel = LEFT;
      WHEN STAGE2 =>
        M3_sel = RIGHT;
    END CASE;
END PROCESS;-- ctrlOut
  
END; 
      
      
